module tb;
    reg clk = 0;
    reg rst = 1;
    wire halted;
    wire [7:0] pc;

    // instanciació del CPU
    cpu uut(.clk(clk), .rst(rst), .halted(halted), .pc_out(pc));

    // toggling clock
    always #5 clk = ~clk; // period 10 time units

    initial begin
        $dumpfile("cpu.vcd");
        $dumpvars(0, tb);
        #12 rst = 0; // treiem reset
        // Fem simulació durant un nombre limitat de cicles
        #1000;
        $finish;
    end
endmodule
